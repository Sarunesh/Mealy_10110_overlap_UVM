`include "uvm_pkg.sv"
import uvm_pkg::*;
`include "mealy_overlap_10110.v"
`include "mealy_overlap_10110_common.sv"
`include "mealy_overlap_10110_intf.sv"
`include "mealy_overlap_10110_tx.sv"
`include "mealy_overlap_10110_seq_lib.sv"
`include "mealy_overlap_10110_sqr.sv"
`include "mealy_overlap_10110_drv.sv"
`include "mealy_overlap_10110_mon.sv"
`include "mealy_overlap_10110_sub.sv"
`include "mealy_overlap_10110_agent.sv"
`include "mealy_overlap_10110_sbd.sv"
`include "mealy_overlap_10110_env.sv"
`include "test_lib.sv"
`include "top.sv"
