interface mealy_overlap_10110_intf(input bit clk, input bit rst);
	logic data_out;
	logic data_in;
endinterface
